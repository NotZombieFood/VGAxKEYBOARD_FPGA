module print(
input [9:0] x, y,
input vidon,
input clk,
input [511:0] mem,
input r, g, b,           /////back_ground
output [9:0] rd_address_mem,
output logic [7:0] red, green, blue 
);

logic [7:0] c_red, c_blue, c_green;
logic p_active;
logic [6:0] linea;
logic [9:0] columna;
logic [7:0] b_red, b_blue, b_green;

 /////////////////Linea//////////////////////////////////////////////////////////////////////////
always_comb begin
	if ( (y >= 31) & ( y < 63) )begin    //Primera linea
		linea = 1;
	end
	else if ( (y >=63) & (y<95)) begin    //segunda linea
		linea = 2;
	end
	else if ( (y >=95) & (y<127)) begin    //Tercera linea
		linea = 3;
	end
	else if ( (y >= 127) &  (y<=159)) begin   //Cuarta linea
		linea = 4;
	end
	else if ( (y >= 159) & (y<191)) begin   //Quinta
		linea = 5;
	end
	else if ( (y >= 191) & (y<223)) begin  //sexta
		linea = 6;
	end
	else if ( (y >= 223) & (y<255)) begin //septima
		linea = 7;
	end
	else if ( (y >= 255) & (y<287)) begin //octava
		linea = 8;
	end
	else if ( (y >= 287) & (y<319)) begin //novena
		linea = 9;
	end
	else if ( (y >= 319) & (y<351)) begin //decima
		linea = 10;
	end
	else if ( (y >= 351) & (y<383)) begin //11
		linea = 11;
	end
	else if ( (y >= 383)& (y<415)) begin //12
		linea = 12;
	end
	else if ( (y >= 415) & (y<447)) begin //13
		linea = 13;
	end
	else if ( (y >= 447)& (y<479)) begin //14
		linea = 14;
	end
	else if ( (y >= 479) & (y<511)) begin //15
		linea = 15;
	end
	else //ninguna
		linea = 0;
end

///////////////////Color de linea/////////////////////////////////////////////////////////
always_comb begin
case (linea)
	1: begin
		c_red = 255;
		c_blue = 0;
		c_green = 0;
	end
	2: begin
		c_red = 0;
		c_blue = 255;
		c_green = 0;
	end
	3: begin
		c_red = 0;
		c_blue = 0;
		c_green = 255;
	end
	4: begin
		c_red = 255;
		c_blue = 255;
		c_green = 0;
	end
	5: begin
		c_red = 255;
		c_blue = 0;
		c_green = 255;
	end
	6: begin
		c_red = 0;
		c_blue = 255;
		c_green = 255;
	end
	7: begin
		c_red = 255;
		c_blue = 255;
		c_green = 255;
	end
	8: begin
		c_red = 120;
		c_blue = 30;
		c_green = 250;
	end
	9: begin
		c_red = 250;
		c_blue = 120;
		c_green = 30;
	end
	10: begin
		c_red = 30;
		c_blue = 250;
		c_green = 120;
	end
	11: begin
		c_red = 89;
		c_blue = 46;
		c_green = 27;
	end
	12: begin
		c_red = 27;
		c_blue = 89;
		c_green = 46;
	end
	13: begin
		c_red = 46;
		c_blue = 27;
		c_green = 89;
	end
	14: begin
		c_red = 200;
		c_blue = 100;
		c_green = 0;
	end
	15: begin
		c_red = 0;
		c_blue = 200;
		c_green = 100;
	end
	default: begin
		c_red = 0;
		c_blue = 0;
		c_green = 0;
	end
endcase
end

////////////////////////columna///////////////////////////////////////////////////////////////
always_comb begin
	if ( (x >= 144) & (x < 160) ) 
		columna = 1;
	else if ( (x >= 160) & (x<176))
		columna = 2;
	else if ( (x >= 176) & (x<192))
		columna = 3;
	else if ( (x >= 192)& (x<208))
		columna = 4;
	else if ( (x >= 208)& (x<224))
		columna = 5;
	else if ( (x >= 224)& (x<240))
		columna = 6;
	else if ( (x >= 240)& (x<256))
		columna = 7;
	else if ( (x >= 256)& (x<272))
		columna = 8;
	else if ( (x >= 272)& (x<288))
		columna = 9;
	else if ( (x >= 288)& (x<304))
		columna = 10;
	else if ( (x >= 304)& (x<320))
		columna = 11;
	else if ( (x >= 320)& (x<336))
		columna = 12;
	else if ( (x >= 336)& (x<352))
		columna = 13;
	else if ( (x >= 352)& (x<368))
		columna = 14;
	else if ( (x >= 368)& (x<384))
		columna = 15;
	else if ( (x >= 384)& (x<400))
		columna = 16;
	else if ( (x >= 400)& (x<416))
		columna = 17;
	else if ( (x >= 416)& (x<432))
		columna = 18;
	else if ( (x >= 432)& (x<448))
		columna = 19;
	else if ( (x >= 448)& (x<464))
		columna = 20;
	else if ( (x >= 464)& (x<480))
		columna = 21;
	else if ( (x >= 480)& (x<496))
		columna = 22;
	else if ( (x >= 496)& (x<512))
		columna = 23;
	else if ( (x >= 512)& (x<528))
		columna = 24;
	else if ( (x >= 528)& (x<544))
		columna = 25;
	else if ( (x >= 544)& (x<560))
		columna = 26;
	else if ( (x >= 560)& (x<576))
		columna = 27;
	else if ( (x >= 576)& (x<592))
		columna = 28;
	else if ( (x >= 592)& (x<608))
		columna = 29;
	else if ( (x >= 608)& (x<624))
		columna = 30;
	else if ( (x >= 624)& (x<640))
		columna = 31;
	else if ( (x >= 640)& (x<656))
		columna = 32;
	else if ( (x >= 656)& (x<672))
		columna = 33;
	else if ( (x >= 672)& (x<688))
		columna = 34;
	else if ( (x >= 688)& (x<704))
		columna = 35;
	else if ( (x >= 704)& (x<720))
		columna = 36;
	else if ( (x >= 720)& (x<736))
		columna = 37;
	else if ( (x >= 736)& (x<752))
		columna = 38;
	else if ( (x >= 752)& (x<768))
		columna = 39;
	else if ( (x >= 768) & (x<784))
		columna = 40;
	else 
		columna = 0;
end

assign rd_address_mem = ((columna - 1) + ((linea - 1)*40));


////////////////////////Asignacion p_active////////////////////////////////////////////////////
assign p_active = mem [ ((x-144-((columna-1)*16)) +  ((y-31-((linea-1)*32))*16))];


////////////////////////////Back_ground/////////////////////////////////////////////

always_comb begin
		if (r)
			b_red = 255;
		else
			b_red = 0;
		if (b)
			b_blue = 255;
		else
			b_blue = 0;
		if (g)
			b_green = 255;
		else 
			b_green = 0;
	end
////////////////////////Asignacion colores de pixel//////////////////////////////////////////////7
always_comb begin
	if (vidon) begin
		if (p_active) begin
			red = c_red;
			blue = c_blue;
			green = c_green;
		end
		else begin
			red = b_red;
			blue = b_blue;
			green = b_green;
		end
	end
	else begin
		red = 0;
		blue = 0;
		green = 0;
	end
end

endmodule 