module rom_1(
	input clk,
	input rst,
	input [9:0] address,
	output [511:0] data
);
logic [511:0] rf [37:0];

always_ff @ (posedge clk) begin
	if (rst) begin
		rf [0] <= 0;
		rf [1] <= 512'b 00000000000000000000000000000000001110000001110000111000000111000011100000011100001110000001110000111000000111000011100000011100001110000001110000111000000111000011100000011100001110000001110000111000000111000011100000011100001111111111110000111111111111000011100000011100001110000001110000111000000111000011100000011100001110000001110000111000000111000011100000011100001110000001110000111000000111000011100000011100000111000011100000001110011100000000011111100000000000011000000000000000000000000000000000000000;   // A
		rf [2] <= 512'b 00000000000000000000000000000000000011111111110000011000000011000011000000001100011000000000110001100000000011000110000000001100011000000000110001100000000011000110000000001100011000000000110001100000000011000011000000001100000110000000110000001111111111000000111111111100000110000000110000110000000011000110000000001100011000000000110001100000000011000110000000001100011000000000110001100000000011000110000000001100011000000000110000110000000011000001100000001100000011111111110000000000000000000000000000000000;  //B
		rf [3] <= 512'b 00000000000000000000000000000000000111111111100000111000000111000011000000011100000000000001110000000000000111000000000000011100000000000001110000000000000111000000000000011100000000000001110000000000000111000000000000011100000000000001110000000000000111000000000000011100000000000001110000000000000111000000000000011100000000000001110000000000000111000000000000011100000000000001110000000000000111000000000000011100000000000001110000110000000111000011100000011100000111111111100000000000000000000000000000000000;  //C  //Esta mal
		rf [4] <= 512'b 00000000000000000000000000000000000111111111110000111000000111000011000000011100001100000001110000110000000111000011000000011100001100000001110000110000000111000011000000011100001100000001110000110000000111000011000000011100001100000001110000110000000111000011000000011100001100000001110000110000000111000011000000011100001100000001110000110000000111000011000000011100001100000001110000110000000111000011000000011100001100000001110000110000000111000011100000011100000111111111110000000000000000000000000000000000;  //D
		rf [5] <= 512'b 00000000000000000000000000000000001111111111110000111000000111000011100000011100000000000001110000000000000111000000000000011100000000000001110000000000000111000000000000011100000000000001110000000000000111000000000000011100000000000001110000000000000111000011111111111100001111111111110000000000000111000000000000011100000000000001110000000000000111000000000000011100000000000001110000000000000111000000000000011100000000000001110000111000000111000011100000011100001111111111110000000000000000000000000000000000;  //E
		rf [6] <= 512'b 00000000000000000000000000000000000000000001110000000000000111000000000000011100000000000001110000000000000111000000000000011100000000000001110000000000000111000000000000011100000000000001110000000000000111000000000000011100000000000001110000000000000111000011111111111100001111111111110000000000000111000000000000011100000000000001110000000000000111000000000000011100000000000001110000000000000111000000000000011100000000000001110000111000000111000011100000011100001111111111110000000000000000000000000000000000;  //F  
		rf [7] <= 512'b 00000000000000000000000000000000000111111111100000110000000111000011000000011100001100000001110000110000000111000011000000011100001100000001110000110000000111000011000000011100001100000001110000110000000111000011001110011100001111111001110000000000000111000000000000011100000000000001110000000000000111000000000000011100000000000001110000000000000111000000000000011100000000000001110000000000000111000000000000011100001110000001110000111000000111000011100000011100000111111111100000000000000000000000000000000000;  //G  
		rf [8] <= 512'b 00000000000000000000000000000000001110000001110000111000000111000011100000011100001110000001110000111000000111000011100000011100001110000001110000111000000111000011100000011100001110000001110000111000000111000011100000011100001110000001110000111111111111000011111111111100001110000001110000111000000111000011100000011100001110000001110000111000000111000011100000011100001110000001110000111000000111000011100000011100001110000001110000111000000111000011100000011100001110000001110000000000000000000000000000000000; //H
		rf [9] <= 512'b 00000000000000000000000000000000000111111111100000011111111110000000001111000000000000111100000000000011110000000000001111000000000000111100000000000011110000000000001111000000000000111100000000000011110000000000001111000000000000111100000000000011110000000000001111000000000000111100000000000011110000000000001111000000000000111100000000000011110000000000001111000000000000111100000000000011110000000000001111000000000000111100000000000011110000000001111111111000000111111111100000000000000000000000000000000000; //I
		rf [10] <= 512'b 00000000000000000000000000000000000000111111100000000011000011000000001100001100000000110000110000000011000011000000001100001100000000110000110000000011000011000000001100001100000000110000110000000011000011000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000111111111100000000000000000000000000000000000; //J
		rf [11] <= 512'b 00000000000000000000000000000000001110000001110000111000000111000001110000011100000111000001110000001110000111000000111000011100000001110001110000000111000111000000001110011100000000111001110000000001110111000000000111011100000000001111110000000000111111000000000011111100000000001111110000000001110111000000000111011100000000111001110000000011100111000000011100011100000001110001110000001110000111000000111000011100000111000001110000011100000111000011100000011100001110000001110000000000000000000000000000000000; //K
		rf [12] <= 512'b 00000000000000000000000000000000001111111111110000111111111111000000000000011100000000000001110000000000000111000000000000011100000000000001110000000000000111000000000000011100000000000001110000000000000111000000000000011100000000000001110000000000000111000000000000011100000000000001110000000000000111000000000000011100000000000001110000000000000111000000000000011100000000000001110000000000000111000000000000011100000000000001110000000000000111000000000000011100000000000001110000000000000000000000000000000000; //L
		rf [13] <= 512'b 00000000000000000000000000000000011000000000011001100000000001100110000000000110011000000000011001100000000001100110000000000110011000000000011001100000000001100110000000000110011000000000011001100000000001100110000110000110011000111100011001100111111001100110011001100110011001100110011001100110011001100110011001100110011011000011011001101100001101100110110000110110011011000011011001101100001101100110110000110110011011000011011001111000000111100111100000011110011110000001111000000000000000000000000000000000; //M
		rf [14] <= 512'b 00000000000000000000000000000000011111000000011001111100000001100111111000000110011111110000011001101111000001100110011100000110011001111000011001100011100001100110001110000110011000111000011001100001110001100110000111000110011000011100011001100001110001100110000111000110011000011100011001100000111001100110000011100110011000001110011001100000111001100110000001110110011000000111011001100000011101100110000001111110011000000011111001100000001111100110000000011110011000000001111000000000000000000000000000000000; //N
		rf [15] <= 512'b 00000000000000000000000000000000000000111100000000001110011100000001100000011000001100000000110000110000000011000011000000001100001100000000110000110000000011000011000000001100001100000000110000110000000011000011000000001100001100000000110000110000000011000011000000001100001100000000110000110000000011000011000000001100001100000000110000110000000011000011000000001100001100000000110000110000000011000011000000001100001100000000110000110000000011000000111001110000000000111100000000000000000000000000000000000000; //O
		rf [16] <= 512'b 00000000000000000000000000000000000000000001110000000000000111000000000000011100000000000001110000000000000111000000000000011100000000000001110000000000000111000000000000011100000000000001110000000000000111000000000000011100000000000001110000000000000111000011111111111100001111111111110000111000000111000011100000011100001110000001110000111000000111000011100000011100001110000001110000111000000111000011100000011100001110000001110000111000000111000011111111111100000111111111100000000000000000000000000000000000; //P
		rf [17] <= 512'b 00000000000000000011000000000000000110111100000000011110011100000011110000001100001111100000110000110110000011000011011000001100001101100000110000110011000011000011001100001100001100110000110000110001100011000011000110001100001100011000110000110000000011000011000000001100001100000000110000110000000011000011000000001100001100000000110000110000000011000011000000001100001100000000110000110000000011000011000000001100001100000000110000011000000110000000111001110000000000111100000000000000000000000000000000000000; //Q
		rf [18] <= 512'b 00000000000000000000000000000000001111000001110000111100000111000011110000011100001111000001110000111100000111000001111000011100000111100001110000011110000111000000111100011100000011110001110000001111000111000000011110011100000001111001110000000111100111000011111111111100001111111111110000111000000111000011100000011100001110000001110000111000000111000011100000011100001110000001110000111000000111000011100000011100001110000001110000111000000111000011111111111100000111111111100000000000000000000000000000000000; //R
		rf [19] <= 512'b 000000000000000000000000000000000000001111110000000011100011100000011100000111000011100000011100001110000000000000111000000000000001110000000000000111000000000000001110000000000000011100000000000001110000000000000011100000000000000111000000000000011100000000000000111000000000000011100000000000000111000000000000011100000000000000111000000000000011100000000000001110000000000000011100000000000001110000111000000111000011110001111000000001111100000000000000000000000000000000000000; //S
		rf [20] <= 512'b 000000000000000000000000000000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000011111111111100001111111111110000000000000000000000000000000000; //T
		rf [21] <= 512'b 00000000000000000000000000000000000000111100000000001110011100000011000000001100001100000000110000110000000011000011000000001100001100000000110000110000000011000011000000001100001100000000110000110000000011000011000000001100001100000000110000110000000011000011000000001100001100000000110000110000000011000011000000001100001100000000110000110000000011000011000000001100001100000000110000110000000011000011000000001100001100000000110000110000000011000011000000001100001100000000110000000000000000000000000000000000; //U
		rf [22] <= 512'b 00000000000000000000000000000000000000011000000000000001100000000000000110000000000000111100000000000011110000000000001111000000000000111100000000000110011000000000011001100000000001100110000000000110011000000000011001100000000011000011000000001100001100000000110000110000000011000011000000001100001100000001100000011000000110000001100000011000000110000001100000011000000110000001100000110000000011000011000000001100001100000000110000110000000011000011000000001100001100000000110000000000000000000000000000000000; //V
		rf [23] <= 512'b 00000000000000000000000000000000000111100111100000110001100011000011000110001100001100011000110000110001100011000011000110001100001100011000110000110001100011000011000110001100001100011000110000110001100011000011000110001100001100011000110000110001100011000011000110001100001100011000110000110001100011000011000110001100001100011000110000110001100011000011000110001100001100011000110000110001100011000011000110001100001100011000110000110001100011000011000110001100001100011000110000000000000000000000000000000000; //W
		rf [24] <= 512'b 00000000000000000000000000000000001100000000110000110000000011000011000000001100000110000001100000011000000110000001100000011000000011000011000000001100001100000000110000110000000011000011000000000110011000000000011001100000000001100110000000000011110000000000001111000000000001100110000000000110011000000000011001100000000011000011000000001100001100000000110000110000000011000011000000011000000110000001100000011000000110000001100000110000000011000011000000001100001100000000110000000000000000000000000000000000; //X //esta mal
		rf [25] <= 512'b 00000000000000000000000000000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000011110000000000001001000000000001100110000000000110011000000000011001100000000011000011000000001100001100000000110000110000000011000011000000011000000110000001100000011000000110000001100000110000000011000011000000001100001100000000110000000000000000000000000000000000; //Y
		rf [26] <= 512'b 000000000000000000000000000000000011111111111100000000000000110000000000000110000000000000011000000000000011000000000000001100000000000001100000000000000110000000000000110000000000000011000000000000011000000000000001100000000000000110000000000000110000000000000011000000000000011000000000000001100000000000000110000000000000110000000000000011000000000000001100000000000001100000000000000110000000000000011000000000000011000000000000001111111111110000000000000000000000000000000000; //z
		rf [27] <= 512'b 00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001100000000000000110000000000000011100000000000001110000000000000000000000000; // ´
		rf [28] <= 512'b 00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000011111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // -
		rf [29] <= 512'b 00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100001111111111110000000000000000000000000000000000001111111111110000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // =
		rf [30] <= 512'b 00000000000000000000000000000000000000111111110000000011000111000000000000011100000000000001110000000000000111000000000000011100000000000001110000000000000111000000000000011100000000000001110000000000000111000000000000011100000000000001110000000000000111000000000000011100000000000001110000000000000111000000000000011100000000000001110000000000000111000000000000011100000000000001110000000000000111000000000000011100000000000001110000000000000111000000001100011100000000111111110000000000000000000000000000000000; // [
		rf [31] <= 512'b 00000000000000000000000000000000001111111100000000111000110000000011100000000000001110000000000000111000000000000011100000000000001110000000000000111000000000000011100000000000001110000000000000111000000000000011100000000000001110000000000000111000000000000011100000000000001110000000000000111000000000000011100000000000001110000000000000111000000000000011100000000000001110000000000000111000000000000011100000000000001110000000000000111000000000000011100011000000001111111100000000000000000000000000000000000000; // ]
		rf [32] <= 512'b 0000000000000000000000000000000000001100000000000000110000000000000011000000000000001100000000000000011000000000000001100000000000000110000000000000001100000000000000110000000000000011000000000000000110000000000000011000000000000001100000000000000011000000000000001100000000000000110000000000000001100000000000000110000000000000011000000000000000110000000000000110000000000000011000000000000000110000000000000011000000000000001100000000000000011000000000000001100000000000000110000000000000000000000000000000000; // \
		rf [33] <= 512'b 00000000000000000000000000000000000000000110000000000000011000000000000011000000000000001100000000000001110000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000001111000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // ;
		rf [34] <= 512'b 00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001100000000000000110000000000000011100000000000001110000000000000000000000000; // '
		rf [35] <= 512'b 00000000000000000000000000000000000000000110000000000000011000000000000011000000000000001100000000000001110000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // ,
		rf [36] <= 512'b 00000000000000000000000000000000000000011000000000000011110000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // .
	   rf [37] <= 512'b 00000000000000000000000000000000000000000000000000000000001100000000000000110000000000000011000000000000011000000000000001100000000000000110000000000000110000000000000011000000000000001100000000000001100000000000000110000000000000011000000000000011000000000000001100000000000000110000000000000110000000000000011000000000000001100000000000001100000000000000110000000000000011000000000000011000000000000001100000000000000110000000000000110000000000000011000000000000001100000000000000000000000000000000000000000000; // /

	end
end

assign data = rf[address];

endmodule 